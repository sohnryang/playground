module top;
  initial begin
    $display("Hell World!");
    $finish;
  end
endmodule
